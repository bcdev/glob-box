netcdf mapped {
dimensions:
	lon = 5 ;
	lat = 5 ;
variables:
	float lon(lon) ;
		lon:long_name = "longitude" ;
		lon:unit = "degrees_east" ;
	float lat(lat) ;
		lat:long_name = "latitude" ;
		lat:unit = "degrees_north" ;
	float CHL1_value(lat, lon) ;
		CHL1_value:parameter_code = "CHL1" ;
		CHL1_value:parameter = "CHL1" ;
		CHL1_value:long_name = "CHL1" ;
		CHL1_value:_FillValue = -999.f ;
		CHL1_value:units = "mg/m3" ;
	short CHL1_flags(lat, lon) ;
		CHL1_flags:parameter_code = "CHL1" ;
		CHL1_flags:parameter = "CHL1" ;
		CHL1_flags:long_name = "CHL1 flags" ;
		CHL1_flags:_FillValue = 0s ;

// global attributes:
		:Conventions = "CF-1.0" ;
		:site_id = "1" ;
		:site_name = "Site Name" ;
		:site_longitude = 0.00f ;
		:site_latitude = 0.00f;
		:site_row = 2s ;
		:site_col = 2s ;
		:netcdf_version = "3.5.1 of Mar 15 2005 16:28:41 $" ;
		:title = "GlobCOLOUR Mapped Test Image" ;
		:grid_type = "Equirectangular" ;
		:lat_step = 1.0f ;
		:lon_step = 1.0f ;
		:max_north_grid = 2.5f ;
		:max_south_grid = -2.5f ;
		:max_west_grid = -2.5f ;
		:max_east_grid = 2.5f ;
		:start_time = "20061124163411" ;
		:end_time = "20061124163414" ;
		:duration_time = 3 ;
data:

 lon = -2.0, -1.0, 0.0, 1.0, 2.0 ;

 lat = 2.0, 1.0, 0.0, -1.0, -2.0 ;

 CHL1_value =
  0.0,   1.0,  2.0,  3.0, 4.0,
  5.0,     _,    _,  8.0, 9.0,
  10.0, 11.0, 12.0, 13.0, 14.0,
  15.0, 16.0, 17.0, 18.0, 19.0,
  20.0, 21.0, 22.0, 23.0, 24.0 ;

CHL1_flags =
  8196, 8196, 8196, 8196, 8196,
  8196,    2,    6, 8196, 8196,
  8196, 8196, 8196, 8196, 8196,
  8196, 8196, 8196, 8196, 8196,
  8196, 8196, 8196, 8196, 8196 ;
}
